library verilog;
use verilog.vl_types.all;
entity ormodule_testbench is
end ormodule_testbench;
