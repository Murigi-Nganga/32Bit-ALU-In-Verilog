library verilog;
use verilog.vl_types.all;
entity ALU32_testbench is
end ALU32_testbench;
