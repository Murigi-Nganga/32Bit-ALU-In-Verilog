library verilog;
use verilog.vl_types.all;
entity andmodule_testbench is
end andmodule_testbench;
