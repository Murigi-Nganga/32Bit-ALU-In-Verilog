//The XOR Module
module xormodule(result,a,b);

input a,b;
output result;

assign result = a ^ b; 

endmodule
