library verilog;
use verilog.vl_types.all;
entity mux4x1module_testbench is
end mux4x1module_testbench;
