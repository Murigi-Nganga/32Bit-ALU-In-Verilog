library verilog;
use verilog.vl_types.all;
entity ALU1_Bit_testbench is
end ALU1_Bit_testbench;
