library verilog;
use verilog.vl_types.all;
entity notmodule_testbench is
end notmodule_testbench;
