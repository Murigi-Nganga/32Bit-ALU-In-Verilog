//The AND Module
module andmodule(result, a, b);
input a,b;
output result;

assign result = a & b;

endmodule
