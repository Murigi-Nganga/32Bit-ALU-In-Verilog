//The Full Adder Module Testbench

`timescale 1ns/1ps

module full_adder_testbench();
reg a,b,cin;
wire sum, cout;

full_adder dut(.a(a), .b(b), .cin(cin), .sum(sum), .cout(cout));
initial begin
		a =1'b0; b=1'b0; cin=1'b0;
		#0.1;
		a =1'b0; b=1'b0; cin=1'b1;
		#0.1;
		a =1'b0; b=1'b1; cin=1'b0;
		#0.1;
		a =1'b0; b=1'b1; cin=1'b1;
		#0.1;
		a =1'b1; b=1'b0; cin=1'b0;
		#0.1;
		a =1'b1; b=1'b0; cin=1'b1;
		#0.1;
		a =1'b1; b=1'b1; cin=1'b0;
		#0.1;
		a =1'b1; b=1'b1; cin=1'b1;		
		#0.1;
	end
	
initial
	begin
		$monitor("Simulation Time = %g, a =%b, b =%b, cin = %b, sum = %b, cout = %b", $time,a,b,cin,sum,cout);
	end
endmodule