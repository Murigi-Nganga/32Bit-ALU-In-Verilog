//The OR Module
module ormodule(result,a,b);
input a, b;
output result;

assign result = a | b;

endmodule