library verilog;
use verilog.vl_types.all;
entity ALU_Bit_MSB_testbench is
end ALU_Bit_MSB_testbench;
