library verilog;
use verilog.vl_types.all;
entity notmodule is
    port(
        result          : out    vl_logic;
        a               : in     vl_logic
    );
end notmodule;
