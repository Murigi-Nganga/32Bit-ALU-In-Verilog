library verilog;
use verilog.vl_types.all;
entity full_adder_testbench is
end full_adder_testbench;
