library verilog;
use verilog.vl_types.all;
entity xormodule_testbench is
end xormodule_testbench;
