library verilog;
use verilog.vl_types.all;
entity mux2x1module_testbench is
end mux2x1module_testbench;
